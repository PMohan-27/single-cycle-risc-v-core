module cpu_top(
    input  clk,
    input  rst
);

 




endmodule