module instr_mem(
    
);


endmodule