module ALU(
    input  [3:0] AluOp,
    input  [31:0] SrcA, SrcB,
    output ZeroFlag, OverflowFlag, NegativeFlag
    output reg [31:0] result
);


endmodule